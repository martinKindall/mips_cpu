`timescale 1ns / 1ps

module regfile(
    
    );
endmodule
